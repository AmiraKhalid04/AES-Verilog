module cipher();
//TODO B: Design this Module
endmodule

//You may need to modifing ports of the functions you use here
//Just Add the ports only