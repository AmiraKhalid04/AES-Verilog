module Cipher();
//TODO B: Design this Module
endmodule

//You may need to modifing ports of the functions you use here
//Just Add the ports only

module InvCipher();
//TODO C: Design this Module
endmodule

//You may need to modifing ports of the functions you use here
//Just Add the ports only

module KeyExpansion();
//TODO D: Design this Module
endmodule

//You may need to modifing ports of the functions you use here
//Just Add the ports only

