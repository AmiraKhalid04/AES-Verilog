module KeyExpansion();
//TODO D: Design this Module
endmodule

//You may need to modifing ports of the functions you use here
//Just Add the ports only