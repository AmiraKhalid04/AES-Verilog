module Cipher();
//TODO B: Design this Module
endmodule

//You may need to modifing ports of the functions you use here
//Just Add the ports only

module InvCipher(
    input [127:0]in ,
    input [127:0]key ,
    output[127:0]out ); //in is Cipher --out is PlainText
//TODO C: Design this Module
   

endmodule


//You may need to modifing ports of the functions you use here
//Just Add the ports only

module KeyExpansion();
//TODO D: Design this Module
endmodule

//You may need to modifing ports of the functions you use here
//Just Add the ports only

