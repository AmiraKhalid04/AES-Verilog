module AddRoundKey ();
    
endmodule


module MixColumns ();
    
endmodule

module InvMixColumns ();
    
endmodule

module ShiftRows ();
    
endmodule

module InvShiftRows ();
    
endmodule

module SubBytes ();
    
endmodule

module InvSubBytes ();
    
endmodule

module RotWord ();
    
endmodule

module SubWord ();
    
endmodule